library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

PACKAGE TYPE_ESTADO_BCD IS
TYPE ESTADO_BCD IS (BCD_0, 
                    BCD_1,
                    BCD_2,
                    BCD_3,
                    BCD_4,
                    BCD_5,
                    BCD_6,
                    BCD_7,
                    BCD_8,
                    BCD_9,);
END PACKAGE TYPE_ESTADO_BCD;