LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; -- USA TODOS OS ELEMENTOS DA LIB IEEE.STD_LOGIC_1164


-- DECLARACAO DE ENTIDADES
ENTITY MEUCIRCUITO2 IS
	PORT (A,B,C,D,E,F: IN STD_LOGIC;
	      Y: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END MEUCIRCUITO2;

--DECLARACAO DE ARQUITETURA
ARCHITECTURE MEUCIRCUITO2_ARCH OF MEUCIRCUITO2 IS
SIGNAL AUX1: STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL AUX1: STD_LOGIC_VECTOR(0 TO 2);
BEGIN
	AUX1 <= A & B & C;
	AUX2 <= D & E & F;
END MEUCIRCUITO2_ARCH;
