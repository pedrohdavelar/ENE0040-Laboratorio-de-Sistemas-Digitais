-- Experimento 06 - Questão 02
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 12/01/2025

-- Registrador de Deslocamento

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY REGISTRADOR_DESLOCAMENTO_BIDIRECIONAL IS
    PORT (CLK, RST, LOAD, DIR, L, R: IN STD_LOGIC;
          D: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
          Q: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END REGISTRADOR_DESLOCAMENTO_BIDIRECIONAL;

ARCHITECTURE ARC_REGISTRADOR_DESLOCAMENTO_BIDIRECIONAL OF REGISTRADOR_DESLOCAMENTO_BIDIRECIONAL IS

SIGNAL GDA_Q : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";

BEGIN
    PROCESS(CLK)
    BEGIN 
        IF RISING_EDGE(CLK) THEN
            IF RST = '1' THEN GDA_Q <= "0000";
            ELSIF LOAD = '1' THEN GDA_Q <= D;
                ELSE CASE DIR IS
                    WHEN '0' => GDA_Q <= GDA_Q(2) & GDA_Q(1) & GDA_Q(0) & L;
                    WHEN '1' => GDA_Q <= R & GDA_Q(3) & GDA_Q(2) & GDA_Q(1);
                    WHEN OTHERS => NULL;
                END CASE;
            END IF;
        END IF;
    END PROCESS;
    Q <= GDA_Q;
END ARC_REGISTRADOR_DESLOCAMENTO_BIDIRECIONAL;     