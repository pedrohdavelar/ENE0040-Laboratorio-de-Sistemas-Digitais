-- Experimento 08 - TESTBENCH Q1
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 05/02/2025

-- Testbench - Tempo de simulação: 310 NS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.TYPE_ESTADO_BCD.ALL;

ENTITY TESTBENCH_E08_BCD_MOD10 IS
END TESTBENCH_E08_BCD_MOD10;

ARCHITECTURE ARC_TESTBENCH_E08_BCD_MOD10 OF TESTBENCH_E08_BCD_MOD10 IS
COMPONENT CONTADOR_BCD_MOD10 IS
    PORT (
        CLOCK   : IN STD_LOGIC;
        RESET   : IN STD_LOGIC;
        ENABLE  : IN STD_LOGIC;
        RCI     : IN STD_LOGIC;
        D       : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        LOAD    : IN STD_LOGIC;
        Q       : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        RCO     : OUT STD_LOGIC;
        CURRENT_STATE: OUT ESTADO_BCD
        );
END COMPONENT;

    SIGNAL CLOCK_TB: STD_LOGIC := '0';
    SIGNAL RESET_TB, ENABLE_TB, RCI_TB, LOAD_TB: STD_LOGIC;
    SIGNAL D_TB: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL Q_TB: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL RCO_TB: STD_LOGIC;
    SIGNAL CURRENT_STATE_TB: ESTADO_BCD;	

    BEGIN
        DUT: CONTADOR_BCD_MOD10 PORT MAP (CLOCK_TB, RESET_TB, ENABLE_TB, RCI_TB, D_TB, LOAD_TB, Q_TB, RCO_TB, CURRENT_STATE_TB);
        CLOCK_TB <= NOT CLOCK_TB AFTER 5 NS;
        PROCESS
        BEGIN
        REPORT "INICIANDO TESTE..." SEVERITY NOTE;
        -- CENARIO 1: CONTAR DE 0 A 9;
        RESET_TB <= '1'; WAIT FOR 10 NS;
        RESET_TB <= '0'; LOAD_TB <= '0'; ENABLE_TB <= '0'; RCI_TB <= '0';
        WAIT FOR 190 NS;
        -- CENARIO 2: LOAD DO NR 5; DEPOIS CONTAR ATE 9
        LOAD_TB <= '1'; D_TB <= "0101"; WAIT FOR 10 NS;
        LOAD_TB <= '0'; WAIT FOR 40 NS;
        -- CENARIO 3: LOAD DO NR 7; DEPOIS ATIVAR RESET PARA SOBRESCREVER O LOAD E DEPOIS CONTAR ATE 9
        LOAD_TB <= '1'; D_TB <= "0111"; WAIT FOR 10 NS;
        RESET_TB <= '1'; WAIT FOR 30 NS;
        LOAD_TB <= '0'; RESET_TB <= '0'; WAIT FOR 20 NS;
        REPORT "TESTE FINALIZADO!" SEVERITY NOTE;
        WAIT;
        END PROCESS;
END ARC_TESTBENCH_E08_BCD_MOD10;