-- Experimento 05 - Questão 01
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 11/12/2024

--SOMADOR DE PALAVRAS DE 4 BITS
--ENTRADA: A E B (4 BITS)
--SAÍDA:       S (5 BITS)

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY E05Q01 IS
	PORT (A,B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	      S:  OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
END E05Q01;

ARCHITECTURE ARC_E05Q01 OF E05Q01 IS
--SOMADOR COMPLETO DO EXPERIMENTO 02 QUESTÃO 01
COMPONENT SOMADOR_COMPLETO is
	PORT (A,B,CIN: IN STD_LOGIC;               --ENTRADAS
      	  S,COUT: OUT STD_LOGIC);                  --SAÍDAS
END COMPONENT;

SIGNAL C1,C2,C3: STD_LOGIC;

BEGIN

SC0: SOMADOR_COMPLETO PORT MAP (A(0),B(0),'0',S(0),C1);
SC1: SOMADOR_COMPLETO PORT MAP (A(1),B(1),C1,S(1),C2);
SC2: SOMADOR_COMPLETO PORT MAP (A(2),B(2),C2,S(2),C3);
SC3: SOMADOR_COMPLETO PORT MAP (A(3),B(3),C3,S(3),S(4));

END ARC_E05Q01;