-- Experimento 04 - Porta OR
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 04/12/2024

-- PORTA OR

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTA_OR IS
	PORT(ENTRADA_1, ENTRADA_2: IN STD_LOGIC;
		 SAIDA_OR:   OUT STD_LOGIC);
END PORTA_OR;

ARCHITECTURE ARC_PORTA_OR OF PORTA_OR IS
BEGIN
	SAIDA_OR <= ENTRADA_1 OR ENTRADA_2;
END ARC_PORTA_OR;