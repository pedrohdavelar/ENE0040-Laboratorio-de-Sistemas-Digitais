-- Experimento 08 - TESTBENCH Q2
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 05/02/2025

-- Testbench - Tempo de simulação: 1110 NS

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.TYPE_ESTADO_BCD.ALL;

ENTITY TESTBENCH_E08_BCD_MOD100 IS
END TESTBENCH_E08_BCD_MOD100;

ARCHITECTURE ARC_TESTBENCH_E08_BCD_MOD100 OF TESTBENCH_E08_BCD_MOD100 IS

COMPONENT CONTADOR_BCD_MOD100 IS
    PORT (
        CLOCK: IN STD_LOGIC;
        RESET: IN STD_LOGIC;
        ENABLE: IN STD_LOGIC;
        D_UNIDADE: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        D_DEZENA: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        LOAD: IN STD_LOGIC;
        Q_UNIDADE: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        Q_DEZENA: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        CURRENT_STATE_UNIDADE: OUT ESTADO_BCD;
        CURRENT_STATE_DEZENA: OUT ESTADO_BCD
        );
END COMPONENT;

SIGNAL CLOCK_TB: STD_LOGIC := '0';
SIGNAL RESET_TB, ENABLE_TB, LOAD_TB: STD_LOGIC;
SIGNAL D_UNIDADE_TB, D_DEZENA_TB: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL Q_UNIDADE_TB, Q_DEZENA_TB: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CURRENT_STATE_UNIDADE_TB, CURRENT_STATE_DEZENA_TB: ESTADO_BCD;

BEGIN
    DUT: CONTADOR_BCD_MOD100 PORT MAP (
        CLOCK_TB, RESET_TB, ENABLE_TB,D_UNIDADE_TB, D_DEZENA_TB,
        LOAD_TB, Q_UNIDADE_TB, Q_DEZENA_TB, CURRENT_STATE_UNIDADE_TB, CURRENT_STATE_DEZENA_TB
    );
    CLOCK_TB <= NOT CLOCK_TB AFTER 5 NS;
    PROCESS
    BEGIN
    REPORT "INICIANDO TESTE..." SEVERITY NOTE;
    -- CENARIO 1: CONTAR DE 0 A 99;
    RESET_TB <= '0'; LOAD_TB <= '0'; ENABLE_TB <= '0';
    WAIT FOR 990 NS;
     -- CENARIO 2: LOAD DOS NUMEROS 19, 28, 37, 46, 55, 64, 73, 82, 91
     RESET_TB <= '0'; LOAD_TB <= '1';
     D_DEZENA_TB <= "0001"; D_UNIDADE_TB <= "1001"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0010"; D_UNIDADE_TB <= "1000"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0011"; D_UNIDADE_TB <= "0111"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0100"; D_UNIDADE_TB <= "0110"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0101"; D_UNIDADE_TB <= "0101"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0110"; D_UNIDADE_TB <= "0100"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "0111"; D_UNIDADE_TB <= "0011"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "1000"; D_UNIDADE_TB <= "0010"; WAIT FOR 10 NS;
     D_DEZENA_TB <= "1001"; D_UNIDADE_TB <= "0001"; WAIT FOR 10 NS;
     -- CENARIO 3: COM A ENTRADA LOAD ATIVA, ATIVAR RESET
     RESET_TB <= '1'; WAIT FOR 30 NS;
    REPORT "TESTE FINALIZADO!" SEVERITY NOTE;
    WAIT;
    END PROCESS;
END ARC_TESTBENCH_E08_BCD_MOD100;