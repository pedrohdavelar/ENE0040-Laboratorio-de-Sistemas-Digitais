-- Experimento 03 - Questão 02
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 13/11/2024

-- Decodificador 4x16
-- Entrada: Vetor A (4bits)
-- Saída: Vetor Y (16 bits)

--Tabela Verdade:
--  A   |          Y
-- 0000    0000 0000 0000 0001  -- 1
-- 0001    0000 0000 0000 0010  -- 2
-- 0010    0000 0000 0000 0100  -- 3
-- 0011    0000 0000 0000 1000  -- 4
-- 0100    0000 0000 0001 0000  -- 5
-- 0101    0000 0000 0010 0000  -- 6
-- 0110    0000 0000 0100 0000  -- 7 
-- 0111    0000 0000 1000 0000  -- 8
-- 1000    0000 0001 0000 0000  -- 9
-- 1001    0000 0010 0000 0000  -- 10
-- 1010    0000 0100 0000 0000  -- 11
-- 1011    0000 1000 0000 0000  -- 12
-- 1100    0001 0000 0000 0000  -- 13
-- 1101    0010 0000 0000 0000  -- 14
-- 1110    0100 0000 0000 0000  -- 15
-- 1111    1000 0000 0000 0000  -- 16


-- Usar atribuições seletivas WITH-SELECT
-- Alterado o nome da entity e da saida Y

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DEC4X16 IS
	PORT (A: IN STD_LOGIC_VECTOR   (3 DOWNTO 0);               -- ENTRADA 4 BITS
      	  Y_DEC: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));          -- SAÍDA 16 BITS
END DEC4X16;

ARCHITECTURE ARC_DEC4X16 OF DEC4X16 IS
BEGIN
    WITH A SELECT
	Y_DEC <= "0000000000000001" WHEN "0000",  -- 1
	         "0000000000000010" WHEN "0001",  -- 2
	         "0000000000000100" WHEN "0010",  -- 3
		     "0000000000001000" WHEN "0011",  -- 4
		     "0000000000010000" WHEN "0100",  -- 5
		     "0000000000100000" WHEN "0101",  -- 6 
		     "0000000001000000" WHEN "0110",  -- 7
		     "0000000010000000" WHEN "0111",  -- 8
		     "0000000100000000" WHEN "1000",  -- 9
		     "0000001000000000" WHEN "1001",  -- 10
		     "0000010000000000" WHEN "1010",  -- 11
		     "0000100000000000" WHEN "1011",  -- 12
		     "0001000000000000" WHEN "1100",  -- 13
		     "0010000000000000" WHEN "1101",  -- 14
		     "0100000000000000" WHEN "1110",  -- 15
		     "1000000000000000" WHEN "1111",  -- 16
		     "0000000000000000" WHEN OTHERS;
END ARC_DEC4X16;