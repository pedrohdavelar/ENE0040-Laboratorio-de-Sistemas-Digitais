-- Experimento 04 - Questão 01
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 27/11/2024

-- Entrada - 3 bits (A,B,C)
-- Saída   - 2 bits (X,Y)

-- X = !ABC + A!B!C + AB
-- Y = !A!B + !AB!C + ABC

-- usar APENAS 2 multiplexadores 4x1 e uma porta inversora

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CIRCUITO_E04Q01 IS
	PORT(A,B,C: IN STD_LOGIC;
		 X,Y:  OUT STD_LOGIC);
END CIRCUITO_E04Q01;

ARCHITECTURE ARC_CIRCUITO_E04Q01 OF CIRCUITO_E04Q01 IS
--Multiplexador 4x1 do Experimento 02 Questão 02
COMPONENT MUX4X1 IS
	PORT (D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);               --ENTRADA
	      S: IN STD_LOGIC_VECTOR (1 DOWNTO 0);               --SELEÇÃO
      	  Y_MUX: OUT STD_LOGIC);
END COMPONENT;	

COMPONENT PORTA_NOT IS
	PORT(ENTRADA: IN STD_LOGIC;
		 SAIDA:   OUT STD_LOGIC);
END COMPONENT;

SIGNAL BARRAMENTOAB: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL BARRAMENTOC_X:  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL BARRAMENTOC_Y:  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL NOT_C: STD_LOGIC;
BEGIN
UX: MUX4X1 PORT MAP(BARRAMENTOC_X,BARRAMENTOAB,X); 
UY: MUX4X1 PORT MAP(BARRAMENTOC_Y,BARRAMENTOAB,Y);
NOT1: PORTA_NOT PORT MAP (C, NOT_C);
BARRAMENTOAB(0) <= B;
BARRAMENTOAB(1) <= A;
BARRAMENTOC_X(0) <= '0';
BARRAMENTOC_X(1) <= C;
BARRAMENTOC_X(2) <= NOT_C;
BARRAMENTOC_X(3) <= '1';
BARRAMENTOC_Y(0) <= '1';
BARRAMENTOC_Y(1) <= NOT_C;
BARRAMENTOC_Y(2) <= '0';
BARRAMENTOC_Y(3) <= C;
END ARC_CIRCUITO_E04Q01;	  