-- Experimento 05 - Questão 02
-- Aluno: Pedro Henrique Dias Avelar 241037112
-- Turma 08
-- Data: 11/12/2024

--SOMADOR DE PALAVRAS DE 4 BITS
--ENTRADA: A E B (4 BITS)
--SAÍDA:       S (5 BITS)

--USAR O OPERADOR '+' DA BIBLIOTECA STD_LOGIC_ARITH

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY E05Q02 IS
	PORT (A,B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	      S:  OUT STD_LOGIC_VECTOR (4 DOWNTO 0));
END E05Q02;

ARCHITECTURE E05Q02_ARC OF E05Q02 IS
BEGIN
S <= ('0' & UNSIGNED(A)) + ('0' & UNSIGNED(B));
END E05Q02_ARC;